`include "addf32.v"

module addf32_tb;
reg[31:0] a,b;
wire[23:0] rm;
wire[31:0] sum;
wire[7:0] l;
addf32 rcaa(a,b,sum);

initial begin
a=0;b=0;
#20 a=32'b01000010101010100100000000000000;b=32'b01000000101000000000000000000000; //+85.125 + 5  = +90.125
#20 a=32'b01000010111111100100000000000000;b=32'b01000000111000000000000000000000; //+127.125 + 7 = +134.125
#20 a=32'b11000001011100100000000000000000;b=32'b11000000101000000000000000000000; //-15.125 - 5  = -20.125
#20 a=32'b01000001011100100000000000000000;b=32'b11000000101000000000000000000000; //+15.125 - 5  = +10.125
#20 a=32'b01000001001100100000000000000000;b=32'b11000000101000000000000000000000; //+11.125 - 5  = +6.125
#20 a=32'b11000001001100100000000000000000;b=32'b01000000101000000000000000000000; //-11.125+5    = -6.125
#20 a=32'b01000001001100100000000000000000;b=32'b01000000101000000000000000000000; //+11.125+5    = +16.125
#20 a=32'b10111111100100000000000000000000;b=32'b11000000101000000000000000000000; //-1.125-5    = -6.125

#20
$finish;

end

initial
$monitor("t=%3d a=%b,b=%b,sum=%b",$time,a,b,sum);

endmodule