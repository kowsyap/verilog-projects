`include "divf32.v"

module divf32_tb;
reg[31:0] a,b;
wire[31:0] div;
wire[23:0] q,r;

divf32 rcaa(a,b,div,q);

initial begin
a=0;b=0;
#20 a=32'b01000010101010100100000000000000;b=32'b01000000101000000000000000000000;  //   85.125 /  5 =  17 
#20 a=32'b01000001011110100000000000000000;b=32'b11000000101000000000000000000000;  //   15.625 / -5 = -3
#20 a=32'b01000001011110100000000000000000;b=32'b01000000101011000000000000000000;  //   15.625 / 5.625 = 2
#20 a=32'b01000000101011000000000000000000;b=32'b01000001011110100000000000000000;  //   5.625 / 15.625 = 0

#20
$finish;

end

initial
$monitor("t=%3d a=%b,b=%b,div=%b,q=%b(%d)",$time,a,b,div,q,q);

endmodule